// seven_segment.v
// Decoder 0..9 -> active-LOW 7-seg (a..g)
module seven_segment (
    input  [3:0] digit,
    output reg [6:0] seg
);

always @(*) begin
    case (digit)
      'b0000 : seg = 7'b1000000;
		'b0001 : seg = 7'b1111001;
		'b0010 : seg = 7'b0100100;
		'b0011 : seg = 7'b0110000;
		'b0100 : seg = 7'b0011001;
		'b0101 : seg = 7'b0010010;
		'b0110 : seg = 7'b0000010;
		'b0111 : seg = 7'b1111000;
		'b1000 : seg = 7'b0000000;
		'b1001 : seg = 7'b0011000;
		'b1010 : seg = 7'b0001000;
		'b1011 : seg = 7'b0000011;
		'b1100 : seg = 7'b1000110;
		'b1101 : seg = 7'b0100001;
		'b1110 : seg = 7'b0000110;
		'b1111 : seg = 7'b0001110;

    endcase
end

endmodule
